*Model Description
.param temp=27


*Including sky130 library files
.lib "sky130_fd_pr/models/sky130.lib.spice" tt


*Netlist Description

XM1 Vdd n1 0 0  sky130_fd_pr__pfet_01v8 w=1 l=0.15

R1 n1 in 55

Vdd vdd 0 -1.8V
Vin  in 0 -1.8V

*simulation commands

.op
.dc Vin 0 -1.8 -0.01

.control

run
display
setplot dc1
.endc

.end

